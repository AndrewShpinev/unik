-------------------------------------------------------------------------------
--
-- Title       : VCC
-- Design      : lab2
-- Author      : user
-- Company     : niiet
--
-------------------------------------------------------------------------------
--
-- File        : c:\Users\student\Desktop\���1\lab2\lab2\src\VCC.vhd
-- Generated   : Fri Feb 10 18:27:52 2017
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {VCC} architecture {VCC}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity VCC is
	 port(
		 Y : out STD_LOGIC
	     );
end VCC;

--}} End of automatically maintained section

architecture VCC of VCC is
begin
	 Y <= ;
	 -- enter your statements here --

end VCC;
